//------------------------------------------------------------------------------
// Copyright 2021 Dominik Salvet
// https://github.com/dominiksalvet/raptorv
//------------------------------------------------------------------------------

module decoder (
    input [31:0] inst
);

endmodule
