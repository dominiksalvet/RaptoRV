// https://github.com/dominiksalvet/RaptoRV

module decoder (
    input [31:0] inst
);

endmodule
