package raptorv_pkg;

    parameter NOP_INST = 32'h13; // todo: check upper zeros

endpackage
