// https://github.com/dominiksalvet/RaptoRV
